LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE pkgTop.ALL;

ENTITY topMOD IS
	PORT(
		indiv0: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		oscraw0: 	INOUT STD_LOGIC;
		oscdiv0: 	INOUT STD_LOGIC;
		CLR: 		IN STD_LOGIC;
		DERECHA:	IN STD_LOGIC;
		IZQUIERDA: 	IN STD_LOGIC;
		CRTL: 		IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DATO:	 	INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		Q: 			INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEG:	 	OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		CD: 		OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE Behavioral OF topMOD IS
BEGIN
	-- OSCILADOR
	OS00:	topdiv00 PORT MAP(
				cdiv0 => indiv0,
				oscout0 => oscraw0,
				outdiv0 => oscdiv0);
	-- REGISTRO UNIVERSAL
	REG0:	Registry PORT MAP(
				CLR => CLR,
				CLK => oscdiv0,
				CD => DERECHA,
				CI => IZQUIERDA,
				CRTL => CRTL,
				DATO => DATO,
				Q => Q);
	
	-- CONVERTIDOR DE BCD A 7 SEGMENTOS
	BCD:	BCD_7SEG PORT MAP(
				BCD => Q,
				SEG => SEG);
END Behavioral;