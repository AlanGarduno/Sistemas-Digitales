LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BIN_MOD IS
    PORT (
        CLK:	 IN  STD_LOGIC;
        CLR:	 IN  STD_LOGIC;
        Y: 		 INOUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		Dato: 	 IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Q: 		 INOUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END ENTITY;
 
ARCHITECTURE Behavioral OF BIN_MOD IS
    -- Se�al temporal para el contador.
    SIGNAL AUX: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
BEGIN
    PROCESS (CLK, CLR, Y) BEGIN
        IF CLR = '0' THEN
            AUX <= "0000";
        ELSIF (CLK'Event and CLK='1')THEN
			IF Y = "00" THEN
				--CONTEO ASCENDENTE
				AUX <= AUX + 1;
			ELSIF Y = "01" THEN
				--CONTEO DESCENDENTE
				AUX <= AUX - 1;
			ELSIF Y = "10" THEN
				--RETENCION DE DATO
				AUX <= Q;
			ELSIF Y = "11" THEN
				--CARGAR DATO
				AUX <= Dato;
			END IF;
        END IF;
    END PROCESS;
 
    Q <= AUX;
END Behavioral;