LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE pkgTop.ALL;
USE packageFF.ALL;

ENTITY topAdder IS
	PORT(
	--	OSCILADOR
		indiv0: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		oscraw0: 	INOUT STD_LOGIC;
		oscdiv0: 	INOUT STD_LOGIC;
	--	REGISTROS
		CLR: 		IN STD_LOGIC;
		DERECHA:	IN STD_LOGIC;
		IZQUIERDA: 	IN STD_LOGIC;
		CRTL: 		IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		A: 			INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		B: 			INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	--	ADDER
		AQ: 		INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		BQ: 		INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		Cf_LED:		INOUT STD_LOGIC;
		S:			INOUT STD_LOGIC;
	--	BCD A 7 SEG
		SQ:			INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEG:	 	OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		CD: 		OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	-- CLR ADDER
		ADD_CLR:	IN STD_LOGIC;
	-- RETENCION DEL REGISTRO SERIAL
		CRTL_S:		IN STD_LOGIC
		);
END ENTITY;

ARCHITECTURE Behavioral OF topAdder IS
-- ENTRADAS Y SALIDAS DEL ADDER
SIGNAL Ci: STD_LOGIC:= '0';
--SIGNAL Cf: STD_LOGIC:= '0'; -- SACAR A UN LED PARA APRECIAR EL DESBORDAMIENTO
-- SE�ALES DEL REGISTRO SERIAL
SIGNAL S_CRTL: STD_LOGIC_VECTOR(1 DOWNTO 0):= "01";	--ROTAR A LA DERECHA
SIGNAL ADD_CLR_CONDITION: STD_LOGIC;
BEGIN
	-- OSCILADOR
	OS00:	topdiv00 PORT MAP(
				cdiv0 => indiv0,
				oscout0 => oscraw0,
				outdiv0 => oscdiv0);
	-- REGISTRO UNIVERSAL
	REGA:	Registry PORT MAP(
				CLR => CLR,
				CLK => oscdiv0,
				CD => DERECHA,
				CI => IZQUIERDA,
				CRTL => CRTL,
				DATO => A,
				Q => AQ);
	-- REGISTRO UNIVERSAL
	REGB:	Registry PORT MAP(
				CLR => CLR,
				CLK => oscdiv0,
				CD => DERECHA,
				CI => IZQUIERDA,
				CRTL => CRTL,
				DATO => B,
				Q => BQ);
	-- FULL ADDER
	ADD0: 	FullAdder PORT MAP(
				A => AQ(0),
				B => BQ(0),
				CLR => ADD_CLR_CONDITION,
				Ci => Ci,
				S => S,
				Cf => Cf_LED);
	--Cf <= Cf_LED;
	-- FLIP FLOP D
	FF_D:	ffD PORT MAP(
				CLR => CLR,
				CLK => oscdiv0,
				D => Cf_LED,
				Q => Ci);
	-- ACARREO
	-- SERIAL REGISTRY
	SREG: 	Registry PORT MAP(
				CLR => ADD_CLR_CONDITION,
				CLK => oscdiv0,
				CD => S,
				CI => OPEN,
				CRTL => S_CRTL,
				DATO => OPEN,
				Q => SQ);
	
	-- CONVERTIDOR DE BCD A 7 SEGMENTOS
	BCD:	BCD_7SEG PORT MAP(
				BCD => SQ,
				SEG => SEG);
	CD <= "1110";
	ADD_CLR_CONDITION<= ADD_CLR OR NOT CRTL(1);
	S_CRTL(0) <= CRTL_S;
END Behavioral;