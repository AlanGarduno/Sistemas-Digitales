LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BIN_GRAY IS
	PORT(
		Q:			IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		G:			INOUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE Behavioral OF BIN_GRAY IS
BEGIN
	--GRAY
		G(3) <= Q(3);
		G(2) <= Q(3) XOR Q(2);
		G(1) <= Q(2) XOR Q(1);
		G(0) <= Q(1) XOR Q(0);
END Behavioral;