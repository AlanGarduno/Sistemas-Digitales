library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity package_dado is

end;

architecture behavioral of package_dado is
begin

end behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity packa_dado is

end;

architecture behavioral of packa_dado is
begin

end behavioral;

