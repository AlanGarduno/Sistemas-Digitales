LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE pkgTop IS
	-- OSCILADOR
	COMPONENT topdiv00 IS
		PORT(
			cdiv0:		IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			oscout0:	INOUT STD_LOGIC;
			outdiv0:	INOUT STD_LOGIC);
	END COMPONENT;
	-- CONVERTIDOR DE BCD A 7 SEGMENTOS
	COMPONENT BCD_7SEG
		PORT(
			BCD:		IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			SEG:		OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;
	-- REGISTRO UNIVERSAL
	COMPONENT Registry IS
		PORT(
			CLR, CLK, CD, CI:	IN STD_LOGIC;
			CRTL:				IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			DATO:				INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Q:					INOUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	-- FULL ADDER
	COMPONENT FullAdder IS
		PORT(
			A,B:	IN STD_LOGIC;
			CLR:	IN STD_LOGIC;
			Ci:		IN STD_LOGIC;
			S,Cf:	OUT STD_LOGIC);
	END COMPONENT;
END pkgTop;